module L2C_normal_loop(


);

endmodule