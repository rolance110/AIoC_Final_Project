module PE_array(

);

endmodule