module L2C_preheat(

);


endmodule