module PPU(



);


endmodule