test 123;
